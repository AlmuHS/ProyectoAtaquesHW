----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    10:59:45 11/22/2020 
-- Design Name: 
-- Module Name:    sistema_clave - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
library UNISIM;
use UNISIM.VComponents.all;

entity sistema_clave is
    Port ( clk : in  STD_LOGIC;
           reset : in  STD_LOGIC;
           req : in  STD_LOGIC;
           data_in : in  STD_LOGIC_VECTOR (3 downto 0);
           ctrl_libre : out  STD_LOGIC;
           ctrl_ok : out  STD_LOGIC;
           ctrl_nok : out  STD_LOGIC;
           ack : out  STD_LOGIC);
end sistema_clave;

architecture Behavioral of sistema_clave is
	component ing_inv_programada is
    Port ( clk : in  STD_LOGIC;
           reset : in  STD_LOGIC;
           req : in  STD_LOGIC;
           clave_in : in  STD_LOGIC_VECTOR (3 downto 0);
           ctrl_libre : out  STD_LOGIC;
           ctrl_ok : out  STD_LOGIC;
           ctrl_nok : out  STD_LOGIC;
           ack : out  STD_LOGIC;
           cont : out  STD_LOGIC_VECTOR (9 downto 0);
           mem : in  STD_LOGIC_VECTOR (3 downto 0));
	end component;

	component ing_inv_cableada is
    Port ( clk : in  STD_LOGIC;
           reset : in  STD_LOGIC;
           req : in  STD_LOGIC;
           data_in : in  STD_LOGIC_VECTOR (3 downto 0);
			  mem	: in std_logic_vector(3 downto 0);
			  --cont_out	: out std_logic_vector(9 downto 0);
			  cont_out	: out std_logic_vector(11 downto 0);
           ctrl_libre : out  STD_LOGIC;
           ctrl_ok : out  STD_LOGIC;
           ctrl_nok : out  STD_LOGIC;
			  ack	: out std_logic);
	end component;
	signal mem			: std_logic_vector(3 downto 0);
	--signal cont_out	: std_logic_vector(9 downto 0);
	signal cont_out	: std_logic_vector(11 downto 0);
	signal cont_out1	: std_logic_vector(11 downto 0);
begin
	ctrl_hw:ing_inv_cableada port map (
		clk => clk,
		reset => reset,
		req => req,
		data_in => data_in,
		mem	=> mem,
		cont_out	=> cont_out,
		ctrl_libre => ctrl_libre,
		ctrl_ok => ctrl_ok,
		ctrl_nok => ctrl_nok,
		ack => ack
	);
--	ctrl_sw:ing_inv_programada port map (
--		clk => clk,
--		reset => reset,
--		req => req,
--		clave_in => data_in,
--		mem	=> mem,
--		cont	=> cont_out,
--		ctrl_libre => ctrl_libre,
--		ctrl_ok => ctrl_ok,
--		ctrl_nok => ctrl_nok,
--		ack => ack
--	);
	
	--cont_out1 <= "00" & cont_out;
	cont_out1 <= cont_out + 1632; --Lee a partir de la posición 32 de la fila 19

	mem_clave:RAMB16_S4
   generic map (
      INIT => X"0", --  Value of output RAM registers at startup
      SRVAL => X"0", --  Output value upon SSR assertion
      WRITE_MODE => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      -- The following INIT_xx declarations specify the initial contents of the RAM
		-- Address 0 to 1023
		INIT_00 => X"9271989923439259073090210044410232768691161862863940366084416071",
		INIT_01 => X"2464136603630834255944909489548453797862649565297565269928814000",
		INIT_02 => X"2752523578908595731727222353612168419537494738056860893468972649",
		INIT_03 => X"7862168224150850064429006590178948556374081237243776281469359725",
		INIT_04 => X"5869533650734488382328140642363533345684095666402885028388444443",
		INIT_05 => X"8017935986540727594154127443649196878879605070234532159769020010",
		INIT_06 => X"5173664004680045880407217910893435250839548305533461176611003175",
		INIT_07 => X"0773160748641008555967031979422447757456277270233323692952118286",
		INIT_08 => X"2076951449793281352198771561046510388375662124905758613483608234",
		INIT_09 => X"4849520466742349341444301024359459420810408487340056212031508424",
		INIT_0A => X"3238057510902863100492023924640886829662410344888716697021901348",
		INIT_0B => X"1034760886991902024910417300042844165835834619724047088177877506",
		INIT_0C => X"9543052503630572906565199471902993572961461644608203877704328338",
		INIT_0D => X"7258762670070537842632204605685616097946383062742066637870027562",
		INIT_0E => X"6541182454635743855376088397555878918654534100863876698527925799",
		INIT_0F => X"2551934941668842997410875705531356291400988992546255499555129929",
		-- Address 1024 to 2047
		INIT_10 => X"9740515873414856035008698393265985910954907145530771363303287626",
		INIT_11 => X"5032773777196404280041913504692000600251596179352280061353944998",
		INIT_12 => X"9923710115497417433639252884861283871156941546494633408586320686",
		INIT_13 => X"4190636368608296306904605286940289711503695231291286555360759767",
		INIT_14 => X"9871363179220868442492372657818339904540417334255045963021047964",
		INIT_15 => X"2270860006591128448627448425542156384044749223451828199293726466",
		INIT_16 => X"1079264603104100863681528348095525501728103348351905547151750012",
		INIT_17 => X"5745103728577917597911692161018552719752907652607134679829486131",
		INIT_18 => X"2697840362738724067731354819265682475743867857074363537462094136",
		INIT_19 => X"1111111111111111111111111115321001111111111111111111111132101210", --selected
		INIT_1A => X"8765615342470312078966446941302283053081336792268655913585264871",
		INIT_1B => X"0281457264291110344065746479559047562424453016760596820423552455",
		INIT_1C => X"9958260039769499020233190885973286633912740866290825986248078262",
		INIT_1D => X"4896422541107140432277510096524676923334951752990223629057771860",
		INIT_1E => X"1841206494182470891183441624051039636264023335274808743805203091",
		INIT_1F => X"5265260136987015266696803657237207986192727957546842791405467997",
		-- Address 2048 to 3071
		INIT_20 => X"2995971306804769046789954624859197843742406829353774356484818665",
		INIT_21 => X"3285143438662834383231712674691820589333332742507403181023572682",
		INIT_22 => X"9808987643116965287125249425837657108609068121518690564151772275",
		INIT_23 => X"3260828424624898488175618812685766263020708458381407070506260608",
		INIT_24 => X"9073725426451747925450016976018809966146553846180066535279194684",
		INIT_25 => X"0336305255663955598983859321065089456231029913214427450960806776",
		INIT_26 => X"7068906893450681817308748299903403794963564525218277160441925790",
		INIT_27 => X"7468751538915303879730107492194606012516568295132522552766535411",
		INIT_28 => X"8973968490058055598395306489774495585467631974382674806756101969",
		INIT_29 => X"5068490366122134557209183850113003198522457323956918567163272322",
		INIT_2A => X"4940435640839909198022784801327321911938063474967419552483856805",
		INIT_2B => X"9119265635566570375153720053136697007962158653330428150008694673",
		INIT_2C => X"4082749739472370847490812724939221781154565019361303127001194218",
		INIT_2D => X"9974268437992117436599284483454935486656003988409077855456077115",
		INIT_2E => X"9591557582929543338288940305600513687761578306351216833444773000",
		INIT_2F => X"1001847131802116186580529549636054319212038026181482814619425365",
		-- Address 3072 to 4095
		INIT_30 => X"5286959066454543326274395171579807304358614892542402115405036666",
		INIT_31 => X"0880818151168174868999992545591866734631330155131456418576401697",
		INIT_32 => X"0905566002934874259966139797837335966239738465554696384103797822",
		INIT_33 => X"2255691347888484343350333163684348515499016846166538690194211736",
		INIT_34 => X"0231130664098896657749908888642468062017570287056506854938784254",
		INIT_35 => X"9960903699945698610190703655091704328311138847050566545432797765",
		INIT_36 => X"4213330993474053159501202897128051057112474133406327198748285721",
		INIT_37 => X"1004030509289547067119873299006400440553295611863823926801470695",
		INIT_38 => X"0428062771454527317696825870740701190208426035642878373853977700",
		INIT_39 => X"7653214973783084204031015313580441666978333022219790506346518692",
		INIT_3A => X"4250987183172275975184553830749738369773567280845084279469176105",
		INIT_3B => X"3523218228341382452679546819091360818119464933057580441503554581",
		INIT_3C => X"9751089282701691409670494862234409163418343676489341304200606331",
		INIT_3D => X"9724613835004941382131631944172620266955955996749524424807052715",
		INIT_3E => X"8322355555895407086321915592569190363044944536770173659037705606",
		INIT_3F => X"1544303104842596899122801713648955928361113182108012037092961556")
   port map (
      DO => mem,      -- 4-bit Data Output
      ADDR => cont_out1,  -- 12-bit Address Input
      CLK => CLK,    -- Clock
      DI => "0000",      -- 4-bit Data Input
      EN => '1',      -- RAM Enable Input
      SSR => reset,    -- Synchronous Set/Reset Input
      WE => '0'       -- Write Enable Input
   );

end Behavioral;

